module MIPS_32Bit (clk);
input clk;
endmodule
