module srg_32Bit_MIPS(clk);
input clk;
endmodule
