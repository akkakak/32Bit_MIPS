module 32Bit_MIPS(clk):

endmodule
